LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE numeric_std.all;

ENTITY circuit IS

PORT();
END circuit;

ARCHITECTURE behaviour OF circuit IS
BEGIN

END behaviour;